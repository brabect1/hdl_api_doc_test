//------------------------------------------------------------
//   Copyright 2010 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

/*
* Class: apb_sequencer
* Sequencer specialization for use with apb_driver.
*
* This implementation is merely a specialization of the default uvm_sequencer
* and would be equally well implemented as a `typedef`.
*/
class apb_sequencer extends uvm_sequencer #(apb_seq_item, apb_seq_item);

// UVM Factory Registration Macro
//
`uvm_component_utils(apb_sequencer)

// Standard UVM Methods:

/*
* Function: new
* Conventional UVM component constructor.
*/
extern function new(string name="apb_sequencer", uvm_component parent = null);

endclass: apb_sequencer

function apb_sequencer::new(string name="apb_sequencer", uvm_component parent = null);
  super.new(name, parent);
endfunction
